module test;
	initial $display("Hello from sysverilog");
endmodule
